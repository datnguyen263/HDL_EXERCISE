library verilog;
use verilog.vl_types.all;
entity d_flipflop_vlg_vec_tst is
end d_flipflop_vlg_vec_tst;
