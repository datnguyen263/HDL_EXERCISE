library verilog;
use verilog.vl_types.all;
entity RAM_IO_vlg_vec_tst is
end RAM_IO_vlg_vec_tst;
