library verilog;
use verilog.vl_types.all;
entity masterslave_dff_vlg_vec_tst is
end masterslave_dff_vlg_vec_tst;
