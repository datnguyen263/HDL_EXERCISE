library verilog;
use verilog.vl_types.all;
entity m21_10bit_vlg_vec_tst is
end m21_10bit_vlg_vec_tst;
