library verilog;
use verilog.vl_types.all;
entity m21 is
    port(
        Y               : out    vl_logic;
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        S               : in     vl_logic
    );
end m21;
