library verilog;
use verilog.vl_types.all;
entity PushdownStack_vlg_vec_tst is
end PushdownStack_vlg_vec_tst;
