library verilog;
use verilog.vl_types.all;
entity dff_setrst_vlg_vec_tst is
end dff_setrst_vlg_vec_tst;
