//module test(sel1, sel0, load, en_ct, D, empty, full, pp, en, reset);
//	input empty, full, pp, en, reset;
//	output sel1, sel0, load, en_ct, D;
//	
//	assign sel1 = ((~empty) & (((~full) & en & (~reset))))
//	assign sel0 =
//	assign load = reset;
//	assign en_ct = 
//	assign D = 
//endmodule
